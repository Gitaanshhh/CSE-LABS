// Simple AND Gate Design
module andGate(x1,x2,f);
input x1, x2;
output f;
and (f, x1, x2);
endmodule
