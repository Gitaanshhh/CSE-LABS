// Q4 (Additional 2)
//x1, x2, x3, and x4, which produces an output value of 1
//whenever three or more of the input variables have the value 1
//IDK YET
module lab4(x1, x2, x3, x4, F);
input x1, x2, x3, x4;
output F;
assign F = (x1 == 0 & )?1:0;
endmodule
